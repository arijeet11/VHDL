library verilog;
use verilog.vl_types.all;
entity gates_vlg_vec_tst is
end gates_vlg_vec_tst;
