LIBRARY ieee;
