library verilog;
use verilog.vl_types.all;
entity gates_vlg_check_tst is
    port(
        c               : in     vl_logic;
        f               : in     vl_logic;
        h               : in     vl_logic;
        k               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end gates_vlg_check_tst;
